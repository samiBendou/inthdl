// Verilog simulation library for c35_IOLIB_ANA_4M
// Owner: austriamicrosystems AG  HIT-Kit: Digital
module APRIO500P (Z,PAD);
  inout Z ;
  inout PAD ;
endmodule
module APRIO50P (Z,PAD);
  inout Z ;
  inout PAD ;
endmodule
module APRIOWP (Z,PAD);
  inout Z ;
  inout PAD ;
endmodule
module AGND3ALLP (VSSA);
  input VSSA ;
endmodule
module AGND5ALLP (VSSA);
  input VSSA ;
endmodule
module AVDD3ALLP (VDDA);
  input VDDA ;
endmodule
module AVDD5ALLP (VDDA);
  input VDDA ;
endmodule
module APRIOP (Z,PAD);
  inout Z ;
  inout PAD ;
endmodule
module APRIO1K5P (Z,PAD);
  inout Z ;
  inout PAD ;
endmodule
module APRIO200P (Z,PAD);
  inout Z ;
  inout PAD ;
endmodule
module ARAILPROT3P;
endmodule
module ARAILPROT5P;
endmodule
